module mod10_counter(rst, clk, count);
    output [3:0] count; //0->9->0
    input clk, rst;
    
    // Code to count
    // and set count back to 0 after 9
endmodule