module mux2to1(m, s, )